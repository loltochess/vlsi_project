module counter_AB cntAB (a_cnt, b_cnt, clk, start);
    output [13-1:0] a_cnt,
    output [8-1:0] b_cnt,
    input clk, start;
    

endmodule
